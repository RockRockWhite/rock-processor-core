// Register with reset value
module REGISTER_R(q, d, rst, clk);
    parameter N = 1;
    parameter INIT = {N{1'b0}};
    output reg [N-1:0] q;
    input [N-1:0]      d;
    input 	      rst, clk;
    initial
        q = INIT;
    always @(posedge clk)
        if (rst)
            q <= INIT;
        else
            q <= d;
endmodule // REGISTER_R
