// Register with reset and clock enable
//  Reset works independently of clock enable
module Register_R_CE (
    q,
    d,
    rst,
    ce,
    clk
);
    parameter N = 1;
    parameter INIT = {N{1'b0}};
    output reg [N-1:0] q;
    input [N-1:0] d;
    input rst, ce, clk;
    initial q = INIT;
    always @(posedge clk)
        if (rst) q <= INIT;
        else if (ce) q <= d;
endmodule  // REGISTER_R_CE
